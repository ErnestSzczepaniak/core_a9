library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity elo is
  port (
  
  );
end entity elo;


architecture rtl of elo is
  
begin
  
  main_proc: process(clk)
  begin
    if rising_edge(clk) then
      if rst = rst_val then
        
      else
        
      end if;
    end if;
  end process main_proc;
  
end architecture rtl;